
module main(
    input logic clk,
    output logic led
);

    blinky blk(clk, led);

endmodule
